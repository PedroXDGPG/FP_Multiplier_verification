interface des_if (input bit clk);
  logic rst;
  logic [7:0] in1;
  logic [7:0] in2;
  logic [8:0] out;
  logic       clk;
endinterface
